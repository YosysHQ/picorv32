`timescale 1 ns / 1 ps
// `define VERBOSE
// `define RANDOM_AXI_DELAYS

module testbench;

	reg clk = 1;
	reg resetn = 0;
	wire trap;

	always #5 clk = ~clk;

	initial begin
		repeat (100) @(posedge clk);
		resetn <= 1;
	end

	wire        mem_axi_awvalid;
	reg         mem_axi_awready = 0;
	wire [31:0] mem_axi_awaddr;
	wire [ 2:0] mem_axi_awprot;

	wire        mem_axi_wvalid;
	reg         mem_axi_wready = 0;
	wire [31:0] mem_axi_wdata;
	wire [ 3:0] mem_axi_wstrb;

	reg  mem_axi_bvalid = 0;
	wire mem_axi_bready;

	wire        mem_axi_arvalid;
	reg         mem_axi_arready = 0;
	wire [31:0] mem_axi_araddr;
	wire [ 2:0] mem_axi_arprot;

	reg         mem_axi_rvalid = 0;
	wire        mem_axi_rready;
	reg  [31:0] mem_axi_rdata;

	picorv32_axi uut (
		.clk            (clk            ),
		.resetn         (resetn         ),
		.trap           (trap           ),
		.mem_axi_awvalid(mem_axi_awvalid),
		.mem_axi_awready(mem_axi_awready),
		.mem_axi_awaddr (mem_axi_awaddr ),
		.mem_axi_awprot (mem_axi_awprot ),
		.mem_axi_wvalid (mem_axi_wvalid ),
		.mem_axi_wready (mem_axi_wready ),
		.mem_axi_wdata  (mem_axi_wdata  ),
		.mem_axi_wstrb  (mem_axi_wstrb  ),
		.mem_axi_bvalid (mem_axi_bvalid ),
		.mem_axi_bready (mem_axi_bready ),
		.mem_axi_arvalid(mem_axi_arvalid),
		.mem_axi_arready(mem_axi_arready),
		.mem_axi_araddr (mem_axi_araddr ),
		.mem_axi_arprot (mem_axi_arprot ),
		.mem_axi_rvalid (mem_axi_rvalid ),
		.mem_axi_rready (mem_axi_rready ),
		.mem_axi_rdata  (mem_axi_rdata  )
	);

	reg [31:0] memory [0:64*1024/4-1];
	initial $readmemh("firmware/firmware.hex", memory);

	reg [63:0] xorshift64_state = 64'd88172645463325252;

	task xorshift64_next;
		begin
			// see page 4 of Marsaglia, George (July 2003). "Xorshift RNGs". Journal of Statistical Software 8 (14).
			xorshift64_state = xorshift64_state ^ (xorshift64_state << 13);
			xorshift64_state = xorshift64_state ^ (xorshift64_state >>  7);
			xorshift64_state = xorshift64_state ^ (xorshift64_state << 17);
		end
	endtask

	reg [2:0] fast_axi_transaction = ~0;
	reg [4:0] delay_axi_transaction = 0;

`ifdef RANDOM_AXI_DELAYS
	always @(posedge clk) begin
		xorshift64_next;
		{fast_axi_transaction, delay_axi_transaction} <= xorshift64_state;
	end
`endif

	reg latched_raddr_en = 0;
	reg latched_waddr_en = 0;
	reg latched_wdata_en = 0;

	reg fast_raddr = 0;
	reg fast_waddr = 0;
	reg fast_wdata = 0;

	reg [31:0] latched_raddr;
	reg [31:0] latched_waddr;
	reg [31:0] latched_wdata;
	reg [ 3:0] latched_wstrb;
	reg        latched_rinsn;

	always @(posedge clk) begin
		mem_axi_arready <= 0;
		mem_axi_awready <= 0;
		mem_axi_wready <= 0;

		fast_raddr <= 0;
		fast_waddr <= 0;
		fast_wdata <= 0;

		if (mem_axi_rvalid && mem_axi_rready) begin
			mem_axi_rvalid <= 0;
		end

		if (mem_axi_bvalid && mem_axi_bready) begin
			mem_axi_bvalid <= 0;
		end

		if (mem_axi_arvalid && mem_axi_arready && !fast_raddr) begin
			latched_raddr = mem_axi_araddr;
			latched_rinsn = mem_axi_arprot[2];
			latched_raddr_en = 1;
		end

		if (mem_axi_awvalid && mem_axi_awready && !fast_waddr) begin
			latched_waddr = mem_axi_awaddr;
			latched_waddr_en = 1;
		end

		if (mem_axi_wvalid && mem_axi_wready && !fast_wdata) begin
			latched_wdata = mem_axi_wdata;
			latched_wstrb = mem_axi_wstrb;
			latched_wdata_en = 1;
		end

		if (mem_axi_arvalid && !(latched_raddr_en || fast_raddr) && !delay_axi_transaction[0]) begin
			mem_axi_arready <= 1;
			if (fast_axi_transaction[0]) begin
				fast_raddr <= 1;
				latched_raddr = mem_axi_araddr;
				latched_rinsn = mem_axi_arprot[2];
				latched_raddr_en = 1;
			end
		end

		if (mem_axi_awvalid && !(latched_waddr_en || fast_waddr) && !delay_axi_transaction[1]) begin
			mem_axi_awready <= 1;
			if (fast_axi_transaction[1]) begin
				fast_waddr <= 1;
				latched_waddr = mem_axi_awaddr;
				latched_waddr_en = 1;
			end
		end

		if (mem_axi_wvalid && !(latched_wdata_en || fast_wdata) && !delay_axi_transaction[2]) begin
			mem_axi_wready <= 1;
			if (fast_axi_transaction[2]) begin
				fast_wdata <= 1;
				latched_wdata = mem_axi_wdata;
				latched_wstrb = mem_axi_wstrb;
				latched_wdata_en = 1;
			end
		end

		if (!mem_axi_rvalid && latched_raddr_en && !delay_axi_transaction[3]) begin
`ifdef VERBOSE
			$display("RD: ADDR=%08x DATA=%08x%s", latched_raddr, memory[latched_raddr >> 2], latched_rinsn ? " INSN" : "");
`endif
			if (latched_raddr < 64*1024) begin
				mem_axi_rdata <= memory[latched_raddr >> 2];
				mem_axi_rvalid <= 1;
				latched_raddr_en = 0;
			end else begin
				$display("OUT-OF-BOUNDS MEMORY READ FROM %08x", latched_raddr);
				$finish;
			end
		end

		if (!mem_axi_bvalid && latched_waddr_en && latched_wdata_en && !delay_axi_transaction[4]) begin
`ifdef VERBOSE
			$display("WR: ADDR=%08x DATA=%08x STRB=%04b", latched_waddr, latched_wdata, latched_wstrb);
`endif
			if (latched_waddr < 64*1024) begin
				if (latched_wstrb[0]) memory[latched_waddr >> 2][ 7: 0] <= latched_wdata[ 7: 0];
				if (latched_wstrb[1]) memory[latched_waddr >> 2][15: 8] <= latched_wdata[15: 8];
				if (latched_wstrb[2]) memory[latched_waddr >> 2][23:16] <= latched_wdata[23:16];
				if (latched_wstrb[3]) memory[latched_waddr >> 2][31:24] <= latched_wdata[31:24];
			end else
			if (latched_waddr == 32'h1000_0000) begin
`ifdef VERBOSE
				if (32 <= latched_wdata && latched_wdata < 128)
					$display("OUT: '%c'", latched_wdata);
				else
					$display("OUT: %3d", latched_wdata);
`else
				$write("%c", latched_wdata);
				$fflush();
`endif
			end else begin
				$display("OUT-OF-BOUNDS MEMORY WRITE TO %08x", latched_waddr);
				$finish;
			end
			mem_axi_bvalid <= 1;
			latched_waddr_en = 0;
			latched_wdata_en = 0;
		end
	end

	initial begin
		$dumpfile("testbench.vcd");
		$dumpvars(0, testbench);
		repeat (1000000) @(posedge clk);
		$display("TIMEOUT");
		$finish;
	end

	always @(posedge clk) begin
		if (resetn && trap) begin
			repeat (10) @(posedge clk);
			$display("TRAP");
			$finish;
		end
	end
endmodule
